*** Figure 1.12 CMOS: Circuit Design, Layout, and Simulation ***

* View listing file to see transfer function information (Edit LL on menu buttons)
.TF 	I(Vmeas) Vin

Vin	Vin	0	DC	1
R1	Vin	Vout	1k
R2	Vout	Vmeas	2k
Vmeas	Vmeas	0	DC	0

.end