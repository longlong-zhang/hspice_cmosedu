*** Figure 1.11_TF CMOS: Circuit Design, Layout, and Simulation ***

* View listing file to see transfer function information (Edit LL on menu buttons)
.TF 	V(Vout,0) 	Vin

Vin	Vin	0	DC	1
R1	Vin	Vout	1k
R2	Vout	0	2k

.end