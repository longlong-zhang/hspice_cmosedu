*** Figure 1.10 CMOS: Circuit Design, Layout, and Simulation ***

* View listing file to see operating point information (Edit LL on menu buttons)
.op

Vin	1	0	DC	1
R1	1	2	1k
R2	2	0	2k

.end